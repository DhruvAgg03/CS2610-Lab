`timescale 1ns/1ns

module MantissaAdder(Sm, Pm, Qm, MAS);

    input[7:0] Pm, Qm;
    input MAS;
    output[8:0] Sm;

    wire[8:0] sum, diff;

    

endmodule