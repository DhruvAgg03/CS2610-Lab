`timescale 1ns/1ns

module ManMul (
    input wire [6:0] Xm, Ym,
    output wire [6:0] Zm,
    output wire PM15
);
    
endmodule