`timescale 1ns/1ns

module ExpAdder (
    input wire [3:0] Xe, Ye,
    input wire PM15,
    output wire [3:0] Ze
);
    
endmodule